module add_1(input [15:0] current, output [15:0] next);
assign next = current + 1'b1;
endmodule
